
interface intf();
    // ------------------- port declaration-------------------------------------
    logic en;
    logic [2:0] in;
    logic [7:0] out;
    //--------------------------------------------------------------------------

endinterface

